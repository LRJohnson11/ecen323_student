package datapathConstants;

    parameter OPCODE_MSB = 6;
    parameter OPCODE_LSB = 0;


endpackage