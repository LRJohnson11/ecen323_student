localparam[3:0] ALUOP_AND = 4'B0000;
localparam[3:0] ALUOP_OR = 4'b0001;
localparam[3:0] ALUOP_ADD = 4'B0010;
localparam[3:0] ALUOP_SUB = 4'b0110;
localparam[3:0] ALUOP_LT = 4'b0111;
localparam[3:0] ALUOP_LSR = 4'b1000;
localparam[3:0] ALUOP_LSL = 4'B1001;
localparam[3:0] ALUOP_ASR = 4'b1010;
localparam[3:0] ALUOP_XOR = 4'b1101;